import rtl_settings_pkg::*;

class statistics;

bit [CSR_RD_REQ : CSR_WR_TICKS][31 : 0] stat_registers;

endclass : statistics
