package tb_settings_pkg;

parameter int CLK_SYS_T = 10_000;
parameter int CLK_MEM_T = 8_000;

parameter int RND_WAITREQ   = 0;
parameter int RND_RVALID    = 0;

parameter int MIN_DELAY_PARAM = 0;
parameter int MAX_DELAY_PARAM = 5;

endpackage : tb_settings_pkg
